`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:57:22 04/05/1612 
// Design Name: 
// Module Name:    display_ctrl 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module display_ctrl(pattern, reset, clk, state);

	input clk;
	input reset;
	input [1:0] state;
	output [255:0] pattern;
	
	reg [255:0] pattern;
	reg [255:0] pattern_next;
	reg [3:0] count;
	reg [3:0] count_next;
	wire [255:0] LG0,LG1,LG2,LG3,LG4,LG5,LG6,LG7,LG8,LG9,LGS;
	
	parameter INIT = 2'b00;
	parameter RUN = 2'b01;
	parameter PAUSE = 2'b10;
	
	always @(posedge clk or negedge reset) begin
		if (reset == 1'b0) begin
			pattern <= 256'd0;
			count <= 4'd0;
		end 
		else begin
			pattern <= pattern_next;
			count <= count_next;
		end
	end
	
	always @(*) begin
		case(state)
			INIT:
				count_next = 0;
			RUN:
				if(count == 4'd10) count_next = 1;
				else count_next = count + 1'b1;
			PAUSE:
				count_next = count;
			default:
				count_next = 0;
		endcase
	end
	
	always @(*) begin
		pattern_next = 256'd0;
		case (count)
			4'd0: pattern_next = LGS;
			4'd1: pattern_next = LG0;
			4'd2: pattern_next = LG1;
			4'd3: pattern_next = LG2;
			4'd4: pattern_next = LG3;
			4'd5: pattern_next = LG4;
			4'd6: pattern_next = LG5;
			4'd7: pattern_next = LG6;
			4'd8: pattern_next = LG7;
			4'd9: pattern_next = LG8;
			4'd10: pattern_next = LG9;
		endcase
	end
	
	assign LG0[15*16+:16] = 16'b0000_0000_0000_0000;
	assign LG0[14*16+:16] = 16'b0000_1100_0000_0000;
	assign LG0[13*16+:16] = 16'b0001_1110_0000_0000;
	assign LG0[12*16+:16] = 16'b0000_1100_0000_0000;
	assign LG0[11*16+:16] = 16'b0000_0110_0000_0000;
	assign LG0[10*16+:16] = 16'b0000_0111_1000_0000;
	assign LG0[ 9*16+:16] = 16'b0000_0111_0100_0000;
	assign LG0[ 8*16+:16] = 16'b0000_1011_0010_0000;
	assign LG0[ 7*16+:16] = 16'b0001_0011_0010_0000;
	assign LG0[ 6*16+:16] = 16'b0000_0011_1000_0000;
	assign LG0[ 5*16+:16] = 16'b0000_0010_1000_0000;
	assign LG0[ 4*16+:16] = 16'b0000_0100_0111_0000;
	assign LG0[ 3*16+:16] = 16'b0000_0100_0000_1000;
	assign LG0[ 2*16+:16] = 16'b0000_0100_0001_0000;
	assign LG0[ 1*16+:16] = 16'b0001_1000_0000_0000;
	assign LG0[ 0*16+:16] = 16'b0000_0000_0000_0000;

	assign LG1[15*16+:16] = 16'b0000_0000_0000_0000;
	assign LG1[14*16+:16] = 16'b0000_1100_0000_0000;
	assign LG1[13*16+:16] = 16'b0001_1110_0000_0000;
	assign LG1[12*16+:16] = 16'b0000_1100_0000_0000;
	assign LG1[11*16+:16] = 16'b0000_0110_0000_0000;
	assign LG1[10*16+:16] = 16'b0000_0111_0000_0000;
	assign LG1[ 9*16+:16] = 16'b0000_0110_1000_0000;
	assign LG1[ 8*16+:16] = 16'b0000_1111_0100_0000;
	assign LG1[ 7*16+:16] = 16'b0001_0011_0100_0000;
	assign LG1[ 6*16+:16] = 16'b0000_0011_1000_0000;
	assign LG1[ 5*16+:16] = 16'b0000_0010_1000_0000;
	assign LG1[ 4*16+:16] = 16'b0000_0100_0110_0000;
	assign LG1[ 3*16+:16] = 16'b0000_1000_0010_0000;
	assign LG1[ 2*16+:16] = 16'b0000_0110_0110_0000;
	assign LG1[ 1*16+:16] = 16'b0000_0010_0000_0000;
	assign LG1[ 0*16+:16] = 16'b0000_1110_0000_0000;

	assign LG2[15*16+:16] = 16'b0000_0000_0000_0000;
	assign LG2[14*16+:16] = 16'b0000_1100_0000_0000;
	assign LG2[13*16+:16] = 16'b0001_1110_0000_0000;
	assign LG2[12*16+:16] = 16'b0000_1100_0000_0000;
	assign LG2[11*16+:16] = 16'b0000_0110_0000_0000;
	assign LG2[10*16+:16] = 16'b0000_0111_0000_0000;
	assign LG2[ 9*16+:16] = 16'b0000_0111_1000_0000;
	assign LG2[ 8*16+:16] = 16'b0000_0111_0100_0000;
	assign LG2[ 7*16+:16] = 16'b0000_0011_0100_0000;
	assign LG2[ 6*16+:16] = 16'b0000_0011_1000_0000;
	assign LG2[ 5*16+:16] = 16'b0000_0010_1000_0000;
	assign LG2[ 4*16+:16] = 16'b0000_0100_0100_0000;
	assign LG2[ 3*16+:16] = 16'b0000_0100_0010_0000;
	assign LG2[ 2*16+:16] = 16'b0000_0100_0001_0000;
	assign LG2[ 1*16+:16] = 16'b0001_1100_0000_1100;
	assign LG2[ 0*16+:16] = 16'b0000_0000_0000_0100;

	assign LG3[15*16+:16] = 16'b0000_0000_0000_0000;
	assign LG3[14*16+:16] = 16'b0000_1100_0000_0000;
	assign LG3[13*16+:16] = 16'b0001_1110_0000_0000;
	assign LG3[12*16+:16] = 16'b0000_1100_0000_0000;
	assign LG3[11*16+:16] = 16'b0000_0110_0000_0000;
	assign LG3[10*16+:16] = 16'b0000_0111_1000_0000;
	assign LG3[ 9*16+:16] = 16'b0000_0111_0100_0000;
	assign LG3[ 8*16+:16] = 16'b0000_1011_0100_0000;
	assign LG3[ 7*16+:16] = 16'b0001_0011_0000_0000;
	assign LG3[ 6*16+:16] = 16'b0000_0011_1000_0000;
	assign LG3[ 5*16+:16] = 16'b0000_0010_1000_0000;
	assign LG3[ 4*16+:16] = 16'b0000_0100_0110_0000;
	assign LG3[ 3*16+:16] = 16'b0000_0100_0001_1000;
	assign LG3[ 2*16+:16] = 16'b0000_0100_0000_1000;
	assign LG3[ 1*16+:16] = 16'b0001_1000_0001_0000;
	assign LG3[ 0*16+:16] = 16'b0000_0000_0000_0000;

	assign LG4[15*16+:16] = 16'b0000_0000_0000_0000;
	assign LG4[14*16+:16] = 16'b0000_1100_0000_0000;
	assign LG4[13*16+:16] = 16'b0001_1110_0000_0000;
	assign LG4[12*16+:16] = 16'b0000_1100_0000_0000;
	assign LG4[11*16+:16] = 16'b0000_0110_0000_0000;
	assign LG4[10*16+:16] = 16'b0000_0111_0000_0000;
	assign LG4[ 9*16+:16] = 16'b0000_0111_0000_0000;
	assign LG4[ 8*16+:16] = 16'b0000_0111_0000_0000;
	assign LG4[ 7*16+:16] = 16'b0000_0011_0000_0000;
	assign LG4[ 6*16+:16] = 16'b0000_0011_0000_0000;
	assign LG4[ 5*16+:16] = 16'b0000_0011_0000_0000;
	assign LG4[ 4*16+:16] = 16'b0000_0011_0000_0000;
	assign LG4[ 3*16+:16] = 16'b0000_0001_0000_0000;
	assign LG4[ 2*16+:16] = 16'b0000_0001_0000_0000;
	assign LG4[ 1*16+:16] = 16'b0000_0001_0000_0000;
	assign LG4[ 0*16+:16] = 16'b0000_0011_0000_0000;

	assign LG5[15*16+:16] = 16'b0000_0000_0000_0000;
	assign LG5[14*16+:16] = 16'b0000_1100_0000_0000;
	assign LG5[13*16+:16] = 16'b0001_1110_0000_0000;
	assign LG5[12*16+:16] = 16'b0000_1100_0000_0000;
	assign LG5[11*16+:16] = 16'b0000_0110_0000_0000;
	assign LG5[10*16+:16] = 16'b0000_0111_1000_0000;
	assign LG5[ 9*16+:16] = 16'b0000_0111_0100_0000;
	assign LG5[ 8*16+:16] = 16'b0000_0111_0010_0000;
	assign LG5[ 7*16+:16] = 16'b0000_1011_0000_0000;
	assign LG5[ 6*16+:16] = 16'b0000_0011_1000_0000;
	assign LG5[ 5*16+:16] = 16'b0000_0010_1000_0000;
	assign LG5[ 4*16+:16] = 16'b0000_0100_0111_0000;
	assign LG5[ 3*16+:16] = 16'b0000_0100_0000_1000;
	assign LG5[ 2*16+:16] = 16'b0001_1100_0000_0000;
	assign LG5[ 1*16+:16] = 16'b0000_0000_0000_0000;
	assign LG5[ 0*16+:16] = 16'b0000_0000_0000_0000;

	assign LG6[15*16+:16] = 16'b0000_0000_0000_0000;
	assign LG6[14*16+:16] = 16'b0000_1100_0000_0000;
	assign LG6[13*16+:16] = 16'b0001_1110_0000_0000;
	assign LG6[12*16+:16] = 16'b0000_1100_0000_0000;
	assign LG6[11*16+:16] = 16'b0000_0110_0000_0000;
	assign LG6[10*16+:16] = 16'b0000_0111_0000_0000;
	assign LG6[ 9*16+:16] = 16'b0000_0110_1000_0000;
	assign LG6[ 8*16+:16] = 16'b0000_0111_1000_0000;
	assign LG6[ 7*16+:16] = 16'b0000_0011_1000_0000;
	assign LG6[ 6*16+:16] = 16'b0000_0011_0000_0000;
	assign LG6[ 5*16+:16] = 16'b0000_0011_0000_0000;
	assign LG6[ 4*16+:16] = 16'b0000_0111_0000_0000;
	assign LG6[ 3*16+:16] = 16'b0000_0100_1000_0000;
	assign LG6[ 2*16+:16] = 16'b0000_0010_0100_0000;
	assign LG6[ 1*16+:16] = 16'b0000_1110_0010_0000;
	assign LG6[ 0*16+:16] = 16'b0000_0000_0000_0000;

	assign LG7[15*16+:16] = 16'b0000_0000_0000_0000;
	assign LG7[14*16+:16] = 16'b0000_1100_0000_0000;
	assign LG7[13*16+:16] = 16'b0001_1110_0000_0000;
	assign LG7[12*16+:16] = 16'b0000_1100_0000_0000;
	assign LG7[11*16+:16] = 16'b0000_0110_0000_0000;
	assign LG7[10*16+:16] = 16'b0000_0111_1000_0000;
	assign LG7[ 9*16+:16] = 16'b0000_0111_0100_0000;
	assign LG7[ 8*16+:16] = 16'b0000_1011_0010_0000;
	assign LG7[ 7*16+:16] = 16'b0001_0011_0010_0000;
	assign LG7[ 6*16+:16] = 16'b0000_0011_1000_0000;
	assign LG7[ 5*16+:16] = 16'b0000_0010_1000_0000;
	assign LG7[ 4*16+:16] = 16'b0000_0100_0110_0000;
	assign LG7[ 3*16+:16] = 16'b0000_0100_0011_0000;
	assign LG7[ 2*16+:16] = 16'b0000_0100_0001_0000;
	assign LG7[ 1*16+:16] = 16'b0001_1000_0010_0000;
	assign LG7[ 0*16+:16] = 16'b0000_0000_0000_0000;

	assign LG8[15*16+:16] = 16'b0000_0000_0000_0000;
	assign LG8[14*16+:16] = 16'b0000_1100_0000_0000;
	assign LG8[13*16+:16] = 16'b0001_1110_0000_0000;
	assign LG8[12*16+:16] = 16'b0000_1100_0000_0000;
	assign LG8[11*16+:16] = 16'b0000_0110_0000_0000;
	assign LG8[10*16+:16] = 16'b0000_0111_0000_0000;
	assign LG8[ 9*16+:16] = 16'b0000_0110_1000_0000;
	assign LG8[ 8*16+:16] = 16'b0000_1111_0100_0000;
	assign LG8[ 7*16+:16] = 16'b0001_0011_0100_0000;
	assign LG8[ 6*16+:16] = 16'b0000_0011_1000_0000;
	assign LG8[ 5*16+:16] = 16'b0000_0010_1000_0000;
	assign LG8[ 4*16+:16] = 16'b0000_0100_0100_0000;
	assign LG8[ 3*16+:16] = 16'b0000_1000_0010_0000;
	assign LG8[ 2*16+:16] = 16'b0000_0110_0001_0000;
	assign LG8[ 1*16+:16] = 16'b0000_0010_0011_0000;
	assign LG8[ 0*16+:16] = 16'b0000_0110_0000_0000;

	assign LG9[15*16+:16] = 16'b0000_0000_0000_0000;
	assign LG9[14*16+:16] = 16'b0000_1100_0000_0000;
	assign LG9[13*16+:16] = 16'b0001_1110_0000_0000;
	assign LG9[12*16+:16] = 16'b0000_1100_0000_0000;
	assign LG9[11*16+:16] = 16'b0000_0110_0000_0000;
	assign LG9[10*16+:16] = 16'b0000_0111_1000_0000;
	assign LG9[ 9*16+:16] = 16'b0000_0111_0100_0000;
	assign LG9[ 8*16+:16] = 16'b0000_1011_0010_0000;
	assign LG9[ 7*16+:16] = 16'b0001_0011_0010_0000;
	assign LG9[ 6*16+:16] = 16'b0000_0011_1000_0000;
	assign LG9[ 5*16+:16] = 16'b0000_0010_1000_0000;
	assign LG9[ 4*16+:16] = 16'b0000_0100_0111_0000;
	assign LG9[ 3*16+:16] = 16'b0000_0100_0000_1000;
	assign LG9[ 2*16+:16] = 16'b0000_0100_0001_0000;
	assign LG9[ 1*16+:16] = 16'b0001_1000_0000_0000;
	assign LG9[ 0*16+:16] = 16'b0000_0000_0000_0000;

	assign LGS[15*16+:16] = 16'b0000_0011_1000_0000;
	assign LGS[14*16+:16] = 16'b0000_0011_1000_0000;
	assign LGS[13*16+:16] = 16'b0000_0011_1000_0000;
	assign LGS[12*16+:16] = 16'b0000_0010_1000_0000;
	assign LGS[11*16+:16] = 16'b0000_0111_1100_0000;
	assign LGS[10*16+:16] = 16'b0000_1111_1110_0000;
	assign LGS[ 9*16+:16] = 16'b0001_1111_1111_0000;
	assign LGS[ 8*16+:16] = 16'b0001_1011_1011_0000;
	assign LGS[ 7*16+:16] = 16'b0001_1011_1011_0000;
	assign LGS[ 6*16+:16] = 16'b0001_1011_1011_0000;
	assign LGS[ 5*16+:16] = 16'b0001_0111_1101_0000;
	assign LGS[ 4*16+:16] = 16'b0000_0110_1100_0000;
	assign LGS[ 3*16+:16] = 16'b0000_0110_1100_0000;
	assign LGS[ 2*16+:16] = 16'b0000_0110_1100_0000;
	assign LGS[ 1*16+:16] = 16'b0000_1110_1110_0000;
	assign LGS[ 0*16+:16] = 16'b0001_1110_1111_0000;
	
	

endmodule












